** Profile: "SCHEMATIC1-bias"  [ C:\Users\Bertan\Desktop\o.c\bias-SCHEMATIC1-bias.sim ] 

** Creating circuit file "bias-SCHEMATIC1-bias.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "D:\DERSLER\5.YARIYIL\EEM 311 LAB\deney 4\deney4\jfet.lib" 
.lib "D:\DERSLER\5.YARIYIL\EEM 311 LAB\deney 3\deney3\cd4007.lib" 
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\bias-SCHEMATIC1.net" 


.END
