** Profile: "SCHEMATIC1-bias"  [ C:\Users\Bertan\Desktop\�.�. 7\oc-schematic1-bias.sim ] 

** Creating circuit file "oc-schematic1-bias.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Windows\pspice.ini file:
.lib "C:\Program Files\OrcadLite\Capture\Library\PSpice\eval.lib" 
.lib "D:\DERSLER\5.YARIYIL\EEM 311 LAB Elektronik II\deney 4\deney4\jfet.lib" 
.lib "D:\DERSLER\5.YARIYIL\EEM 311 LAB Elektronik II\deney 3\deney3\cd4007.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\oc-SCHEMATIC1.net" 


.END
