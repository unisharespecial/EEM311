** Profile: "SCHEMATIC1-deney3"  [ C:\Documents and Settings\MR.ERAY\Desktop\EEM311- ELEKTRONIK 2\LABS\deney3\deney3-schematic1-deney3.sim ] 

** Creating circuit file "deney3-schematic1-deney3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of pspiceev.ini file:
.lib "C:\Documents and Settings\MR.ERAY\Desktop\EEM311- ELEKTRONIK 2\LABS\deney3\cd4007.lib" 
.lib "C:\Documents and Settings\MR.ERAY\Desktop\EEM311- ELEKTRONIK 2\LABS\deney1\deney1\EEM311.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 15ms 0 10us 
.PROBE 
.INC "deney3-SCHEMATIC1.net" 

.INC "deney3-SCHEMATIC1.als"


.END
