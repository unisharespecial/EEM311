** Profile: "SCHEMATIC1-sim1"  [ C:\Documents and Settings\LuCiFeR\Desktop\deney6 pspice\aaaaaaa-schematic1-sim1.sim ] 

** Creating circuit file "aaaaaaa-schematic1-sim1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "C:\Documents and Settings\LuCiFeR\Desktop\deney6\cd4007.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3ms 0 1uF 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\aaaaaaa-SCHEMATIC1.net" 


.END
