** Profile: "SCHEMATIC1-deney7"  [ C:\Documents and Settings\Tolga Aydin\Desktop\eem311fb\deney7-schematic1-deney7.sim ] 

** Creating circuit file "deney7-schematic1-deney7.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "C:\Documents and Settings\Tolga Aydin\Desktop\deney4\jfet.lib" 
.lib "C:\Documents and Settings\Tolga Aydin\Desktop\deney6\cd4007.lib" 
.lib "C:\Documents and Settings\Tolga Aydin\Desktop\deney1\EEM311.lib" 
.lib "C:\Program Files\OrcadLite\Capture\Library\PSpice\diode.lib" 
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\deney7-SCHEMATIC1.net" 


.END
